module MMC1 (
    map_bus.mapper bus
);

endmodule
