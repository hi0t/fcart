module chr_ram #(
    parameter ADDR_BITS = 23  // SDRAM width + 1
) (
    input logic clk,
    input logic reset,
    sdram_bus.controller ram,

    input logic [ADDR_BITS-1:0] addr,
    input logic [7:0] data_in,
    output logic [7:0] data_out,
    input logic ce,
    input logic oe,
    input logic we
);
    logic [1:0] read_sync;
    logic [3:0] write_sync;
    logic [2:0][ADDR_BITS-1:0] addr_gray;
    logic [2:0] match_addr;

    assign data_out = addr[0] ? ram.data_read[15:8] : ram.data_read[7:0];

    always_ff @(posedge clk) begin
        if (reset) begin
            ram.req <= 0;
            ram.we <= 0;
            read_sync <= '0;
            write_sync <= '0;
            addr_gray <= '1;
            match_addr <= '0;
        end else begin
            read_sync  <= {read_sync[0], ce && !oe};
            write_sync <= {write_sync[2:0], ce && we};
            addr_gray  <= {addr_gray[1:0], addr ^ (addr >> 1)};

            if (read_sync[1] && addr_gray[2] == addr_gray[1]) begin
                match_addr <= {match_addr[1:0], 1'b1};
            end else begin
                match_addr <= '0;
            end

            if (ram.req == ram.ack && match_addr == 3'b011) begin
                ram.we <= 0;
                ram.address <= addr[ADDR_BITS-1:1];
                ram.req <= !ram.req;
            end else if (ram.req == ram.ack && write_sync[3:1] == 3'b100) begin
                ram.we <= 1;
                ram.address <= addr[ADDR_BITS-1:1];
                ram.data_write <= {data_in, data_in};
                ram.wm <= addr[0] ? 2'b01 : 2'b10;
                ram.req <= !ram.req;
            end
        end
    end

`ifdef DEBUG
    logic debug_ram_busy = ram.req != ram.ack;
    logic debug_ram_we = ram.we;
`endif
endmodule
