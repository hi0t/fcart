// GSR blackbox
// verilator lint_off UNUSEDSIGNAL
// verilator lint_off UNDRIVEN

module GSR (GSR);
    input GSR;
endmodule
