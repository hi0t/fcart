// PLL blackbox
// verilator lint_off UNUSEDSIGNAL
// verilator lint_off UNDRIVEN

module pll (inclk0, c0, locked);
    input inclk0;
    output c0;
    output locked;
endmodule
