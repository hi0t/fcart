module fcart (
    input  logic CLK_IN,
    output logic FPGA_IRQ,

    // QSPI
    input logic QSPI_CLK,
    input logic QSPI_NCS,
    inout wire [3:0] QSPI_IO,

    // SDRAM
    output logic SDRAM_CLK,
    output logic SDRAM_CS,
    output logic [11:0] SDRAM_ADDR,
    output logic [1:0] SDRAM_BA,
    inout wire [15:0] SDRAM_DQ,
    output logic SDRAM_RAS,
    output logic SDRAM_CAS,
    output logic SDRAM_WE,
    output logic [1:0] SDRAM_DQM,

    // Cart
    input logic M2,
    input logic [14:0] CPU_ADDR,
    inout wire [7:0] CPU_DATA,
    input logic CPU_RW,
    input logic ROMSEL,
    output logic IRQ,
    input logic PPU_RD,
    input logic PPU_WR,
    output logic CIRAM_A10,
    output logic CIRAM_CE,
    input logic [13:0] PPU_ADDR,
    inout wire [7:0] PPU_DATA,
    output logic SND_OUT,
    output logic CPU_DIR,
    output logic PPU_DIR
);
    localparam RAM_ADDR_BITS = 22;  // SDRAM row + col + bank bits

    logic clk;
    logic async_nreset;
    logic reset;
    logic [7:0] cpu_data_out;
    logic [7:0] ppu_data_out;
    logic [31:0] wr_reg;
    logic [3:0] wr_reg_addr;
    logic wr_reg_changed;
    logic [31:0] launcher_status;
    logic sdram_refresh;
    logic [15:0] pcm;
    logic [7:0] joy1;

    assign CPU_DATA = CPU_DIR ? cpu_data_out : 'z;
    assign PPU_DATA = PPU_DIR ? ppu_data_out : 'z;

    joy_snoop joy (
        .m2(M2),
        .cpu_addr({!ROMSEL, CPU_ADDR}),
        .cpu_data(CPU_DATA[0]),
        .cpu_rw(CPU_RW),
        .joy1(joy1)
    );

    sdram_bus #(.ADDR_BITS(RAM_ADDR_BITS)) ch_ppu (), ch_cpu (), ch_api ();

    map_mux mux (
        .clk(clk),
        .ch_prg(ch_cpu.controller),
        .ch_chr(ch_ppu.controller),
        .refresh(sdram_refresh),

        .m2(M2),
        .cpu_addr({!ROMSEL, CPU_ADDR}),
        .cpu_data_in(CPU_DATA),
        .cpu_data_out(cpu_data_out),
        .cpu_rw(CPU_RW),
        .irq(IRQ),
        .ppu_rd(PPU_RD),
        .ppu_wr(PPU_WR),
        .ciram_a10(CIRAM_A10),
        .ciram_ce(CIRAM_CE),
        .ppu_addr(PPU_ADDR),
        .ppu_data_in(PPU_DATA),
        .ppu_data_out(ppu_data_out),

        .cpu_dir(CPU_DIR),
        .ppu_dir(PPU_DIR),

        .wr_reg(wr_reg[14:0]),
        .wr_reg_addr(wr_reg_addr),
        .wr_reg_changed(wr_reg_changed),
        .status_reg(launcher_status),
        .audio(pcm),
        .joy1(joy1)
    );

    snd_dac snd_dac (
        .m2(M2),
        .pcm_in(pcm),
        .volume(8'd255),
        .pdm_out(SND_OUT)
    );

    pll pll (
        .CLKI (CLK_IN),
        .CLKOP(clk),
        .CLKOS(SDRAM_CLK),
        .LOCK (async_nreset)
    );
    logic [1:0] rst_sync;
    assign reset = !rst_sync[1];
    always_ff @(posedge clk) begin
        if (!async_nreset) begin
            rst_sync <= 2'b00;
        end else begin
            rst_sync <= {rst_sync[0], 1'b1};
        end
    end

    sdram sdram (
        .clk(clk),
        .reset(reset),
        .ch0(ch_cpu.memory),
        .ch1(ch_ppu.memory),
        .ch2(ch_api.memory),
        .refresh(sdram_refresh),
        .sdram_cs(SDRAM_CS),
        .sdram_addr(SDRAM_ADDR),
        .sdram_ba(SDRAM_BA),
        .sdram_dq(SDRAM_DQ),
        .sdram_ras(SDRAM_RAS),
        .sdram_cas(SDRAM_CAS),
        .sdram_we(SDRAM_WE),
        .sdram_dqm(SDRAM_DQM)
    );

    logic [15:0] qspi_rd_data;
    logic qspi_rd_valid;
    logic qspi_rd_ready;
    logic [15:0] qspi_wr_data;
    logic qspi_wr_valid;
    logic qspi_wr_ready;
    logic qspi_start;
    qspi qspi (
        .clk(clk),
        .async_reset(!async_nreset),

        .qspi_clk(QSPI_CLK),
        .qspi_ncs(QSPI_NCS),
        .qspi_io (QSPI_IO),

        .rd_data(qspi_rd_data),
        .rd_valid(qspi_rd_valid),
        .rd_ready(qspi_rd_ready),
        .wr_data(qspi_wr_data),
        .wr_valid(qspi_wr_valid),
        .wr_ready(qspi_wr_ready),
        .start(qspi_start)
    );

    api api (
        .clk(clk),
        .reset(reset),
        .fpga_irq(FPGA_IRQ),

        .wr_reg(wr_reg),
        .wr_reg_addr(wr_reg_addr),
        .wr_reg_changed(wr_reg_changed),
        .ev_reg(launcher_status),

        .ram(ch_api.controller),

        .rd_data(qspi_rd_data),
        .rd_valid(qspi_rd_valid),
        .rd_ready(qspi_rd_ready),
        .wr_data(qspi_wr_data),
        .wr_valid(qspi_wr_valid),
        .wr_ready(qspi_wr_ready),
        .start(qspi_start)
    );
endmodule
